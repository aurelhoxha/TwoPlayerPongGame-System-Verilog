`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 12/17/2016 01:06:59 PM
// Design Name: 
// Module Name: JoinerXOX
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


/*module JoinerXOX(
    input logic [1:0] rows, columns, input logic start,
                    input logic clk, output logic shcp, stcp, mr, oe, ds,[7:0] rowsOut
    );
    logic [7:0][23:0] board;
    TwoPlayerJoiner  gameXOX(rows, columns,start, clk,board );
    Gametop lightTheLedsUp(shcp, stcp, mr, oe, ds,rowsOut, clk, board);
endmodule*/
